//4 BIT UP/DOWN COUNTER 
module updowncounter(clk,rst,ud,out); 
input clk,rst,ud; 
output reg[3:0]out = 4’b0000;


endmodule
